module PD(clk, rst_n, data, flag, addr, fin);
    input clk;
    input rst_n;
    input [9:0]data;
    output flag;
    output [9:0]addr;
    output fin;
    //code here
endmodule
