module LPD(clk, rst_n, data, flag, addr, fin, count);
    input clk;
    input rst_n;
    input [9:0]data;
    output flag;
    output [9:0]addr;
    output fin;
    output [3:0]count;
    //your code
endmodule
